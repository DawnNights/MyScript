module ast